`define OPCODE 6:0
`define    